`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:18:13 08/31/2022 
// Design Name: 
// Module Name:    wrapper_cla_4bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module wrapper_cla_4bit(input clk, input rst, input [3:0] in1, input [3:0] in2, input cin, output reg [3:0] sum, output reg cout)

	reg 

endmodule
